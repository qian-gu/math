package math_pkg;

    `define MATH_MULT_USE_MBE_IV;

endpackage
