package math;

endpackage
