package math_pkg;

  // different modified booth encoding
  typedef enum integer {
      MBE_I   = 0,
      MBE_II  = 1,
      MBE_III = 2,
      MBE_IV  = 3
  } mbe_e;

endpackage
